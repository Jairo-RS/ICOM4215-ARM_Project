`include "CPU.v"

module main;

endmodule
